library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity CLK_GEN is
end CLK_GEN;

architecture rtl of CLK_GEN is

begin


end rtl;

